module top_module (
    output out);

    wire out_wire = 1'b0;
    assign out = out_wire;

endmodule
